module stc ();

endmodule // stc
