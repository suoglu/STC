// This module simulates a sea clutter and radar interface
// 50MHz clock freq

module radar(arp, acp, trig, rst, clk)
input clk, rst;
output reg acp, trig;
output arp;



endmodule
