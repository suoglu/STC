// This module simulates a sea clutter and radar interface

